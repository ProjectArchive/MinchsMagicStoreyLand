NETWORK OF RESISTORS AND DEPENDENT SOURCES
*
* Reduce this complicated collection of dependencies
* down to a single Thevenin equivalent between node 2 and
* the ground node 0
*
I1 1 4 2
V1 1 0 5
E1 5 2 1 3 0.4
F1 5 6 R1 3e-2
G1 2 3 4 6 1.3
H1 3 0 R3 1
R1 4 5 2.2
R2 1 2 470
R3 0 2 330
R4 3 6 22k
R5 5 6 1e4
*
* Look at the voltage at node 2 and the impedance looking into node 2
*
.print dc v(2) z(2)
.dc
.end
