DIODE CASCADE

.model 1N414 D IS=2e-14

Vcc 1 0 5
Dx 1 10 1N414
Dy 10 20 1N414
Dz 20 30 1N414
Rd1 10 0 1k
Rd2 20 0 1k
Rd3 30 0 1k

.print dc v(10) v(20) v(30)
.dc Vcc 0 5 0.5 >eg6.dat
.end
