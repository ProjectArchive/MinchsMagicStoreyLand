#RESISTOR DRIVEN BY VOLTAGE SOURCE
Vsupply ( 0 2 )  DC  10.
R1 ( 0 2 )  1000
