#RESISTOR DRIVEN BY VOLTAGE SOURCE
Vsupply ( 0 2 )  DC  10.
Rc ( 0 2 )  1000
