.TITLE Basic RC Circuit

Vin 0 1 AC 1.5
R1 1 2 1K
C1 1 0 1UF

.OPTION OUT=80
.PRINT OP Iter(0) V(1)

.PLOT AC VDB(1)(-20,0)

.AC 5 1K OCT
